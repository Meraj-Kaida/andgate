module andgate(a,b,y);
input a,b;
output y;
  //jjjjjjj
assign y= a&b;
  //made and gate
endmodule
